
`include "uvm_macros.svh"
import uvm_pkg::*;

interface add_if;
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] y;
endinterface
